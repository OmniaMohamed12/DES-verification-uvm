package DES_Package;
    `include"uvm_macros.svh"
    import uvm_pkg::*;
    `include "DES_Seq_Item.svh"
    `include "DES_Sequences.svh"
    `include "DES_Seq_Library.svh"
    `include "DES_Driver.svh"
    `include "DES_Monitor.svh"
    `include "DES_Sequencer.svh"
    `include "DES_Agent_Config.svh"
    `include "DES_Agent.svh"
    `include "DES_Scoreboard.svh"
    `include "DES_Subscriber.svh"
    `include "DES_Env_Config.svh"
    `include "DES_Env.svh"
    `include "DES_Test.svh"
endpackage